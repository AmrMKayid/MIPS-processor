/**
  * The control unit of a MIPS processor 
  * Input: Opcode of the instruction
  * 
  * Nine single-bit singals: 
  * 1) RegDst
  * 2) RegWrite
  * 3) ALUSrc
  * 4) PCsrc
  * 5) MemRead
  * 6) MemWrite
  * 7) MemtoReg
  * 8) ALU op
  * 9) ALU op
  */

module ControlUnit(RegDst, RegWrite, ALUSrc, Branch, MemRead, MemWrite, MemtoReg, ALUop, OPCode);

	output reg RegDst, RegWrite, ALUSrc, Branch, MemRead, MemWrite, MemtoReg;
	output reg[1:0] ALUop;
	input [5:0] OPCode;

	always@(OPCode) begin
		case(OPCode)
		6'h00: RegDst <= 1; RegWrite <= 1; ALUSrc <= 0; Branch <= 0; MemRead <= 0; MemWrite <= 0; MemtoReg <= 0; ALUop <= 2; /*R instructions*/
		6'h08: RegDst <= 0; RegWrite <= 1; ALUSrc <= 1; Branch <= 0; MemRead <= 0; MemWrite <= 0; MemtoReg <= 0; ALUop <= 2; /*Addi*/ 
		6'h23: RegDst <= 0; RegWrite <= 1; ALUSrc <= 1; Branch <= 0; MemRead <= 1; MemWrite <= 0; MemtoReg <= 1; ALUop <= 0; /*lw*/ 
		6'h2B: RegDst <= 0; RegWrite <= 0; ALUSrc <= 1; Branch <= 0; MemRead <= 0; MemWrite <= 1; MemtoReg <= 0; ALUop <= 0; /*sw*/ 
		6'h21: RegDst <= 0; RegWrite <= 1; ALUSrc <= 1; Branch <= 0; MemRead <= 1; MemWrite <= 0; MemtoReg <= 1; ALUop <= 0; /*lh*/ 
		6'h25: RegDst <= 0; RegWrite <= 1; ALUSrc <= 1; Branch <= 0; MemRead <= 1; MemWrite <= 0; MemtoReg <= 1; ALUop <= 0; /*lhu*/
		6'h0C: RegDst <= 0; RegWrite <= 1; ALUSrc <= 1; Branch <= 0; MemRead <= 0; MemWrite <= 0; MemtoReg <= 0; ALUop <= 2; /*andi*/ 
		6'h0D: RegDst <= 0; RegWrite <= 1; ALUSrc <= 1; Branch <= 0; MemRead <= 0; MemWrite <= 0; MemtoReg <= 0; ALUop <= 2; /*ori*/
		6'h04: RegDst <= 0; RegWrite <= 0; ALUSrc <= 0; Branch <= 1; MemRead <= 0; MemWrite <= 0; MemtoReg <= 0; ALUop <= 1; /*beq*/
		endcase

	end


endmodule