/**
  * Processor Module
  *
  * single cycle MIPS processor module 
  *
  */

module Processor();

	wire[32] pc;

	ProgramCounter PC(pc, PrevPC, clk);
	





endmodule